module moduloControladorJuego (reloj, reinicio, botonArriba, botonAbajo, botonIzquierda, botonDerecha, tableroJuego, estadoJuego);
	input logic reloj;
	input logic reinicio;
	input logic botonArriba;
	input logic botonAbajo;
	input logic botonIzquierda;
	input logic botonDerecha;
	output logic [3:0] tableroJuego [3:0][3:0];
	output logic [1:0] estadoJuego;

	reg [2:0] ESTADO_ACTUAL;
	reg [21:0] CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_COLUMNA_ALEATORIA;
	reg [18:0] CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_FILA_ALEATORIA;
	reg [1:0] POSICION_COLUMNA_ALEATORIA;
	reg [1:0] POSICION_FILA_ALEATORIA;
	
	reg [1:0] POSICION_COLUMNA_ANALIZADA;
	reg [1:0] POSICION_FILA_ANALIZADA;

	parameter [3:0] ESTADO_INICIANDO_JUEGO = 4'b0000;
	parameter [3:0] ESTADO_ESPERANDO_MOVIMIENTO = 4'b0001;
	parameter [3:0] ESTADO_MOVIENDO_HACIA_ARRIBA = 4'b0010;
	parameter [3:0] ESTADO_MOVIENDO_HACIA_ABAJO = 4'b0011;
	parameter [3:0] ESTADO_MOVIENDO_HACIA_IZQUIERDA = 4'b0100;
	parameter [3:0] ESTADO_MOVIENDO_HACIA_DERECHA = 4'b0101;
	parameter [3:0] ESTADO_VERIFICANDO_GANAR_PERDER = 4'b0110;
	parameter [3:0] ESTADO_GENERANDO_POSICION_ALEATORIA = 4'b0111;
	parameter [3:0] ESTADO_GANAR = 4'b1000;
	parameter [3:0] ESTADO_PERDER = 4'b1001;

	always @(posedge reloj) begin
		if (reinicio == 1'b1) begin
			tableroJuego[0][0] <= 4'b0000;
			tableroJuego[0][1] <= 4'b0000;
			tableroJuego[0][2] <= 4'b0000;
			tableroJuego[0][3] <= 4'b0000;
			tableroJuego[1][0] <= 4'b0000;
			tableroJuego[1][1] <= 4'b0000;
			tableroJuego[1][2] <= 4'b0000;
			tableroJuego[1][3] <= 4'b0000;
			tableroJuego[2][0] <= 4'b0000;
			tableroJuego[2][1] <= 4'b0000;
			tableroJuego[2][2] <= 4'b0000;
			tableroJuego[2][3] <= 4'b0000;
			tableroJuego[3][0] <= 4'b0000;
			tableroJuego[3][1] <= 4'b0000;
			tableroJuego[3][2] <= 4'b0000;
			tableroJuego[3][3] <= 4'b0000;
			estadoJuego = 2'b00;
			ESTADO_ACTUAL = ESTADO_INICIANDO_JUEGO;
		end
		else begin
			if (ESTADO_ACTUAL == ESTADO_INICIANDO_JUEGO) begin
				tableroJuego[POSICION_FILA_ALEATORIA][POSICION_COLUMNA_ALEATORIA] = 4'b0001;
				ESTADO_ACTUAL = ESTADO_ESPERANDO_MOVIMIENTO;
			end
			
			if (ESTADO_ACTUAL == ESTADO_ESPERANDO_MOVIMIENTO) begin
				if (botonArriba == 1'b1) begin
					ESTADO_ACTUAL <= ESTADO_MOVIENDO_HACIA_ARRIBA;
					POSICION_COLUMNA_ANALIZADA <= 2'b00;
					POSICION_FILA_ANALIZADA <= 2'b11;
				end
				else if (botonAbajo == 1'b1) begin
					ESTADO_ACTUAL <= ESTADO_MOVIENDO_HACIA_ABAJO;
					POSICION_COLUMNA_ANALIZADA <= 2'b00;
					POSICION_FILA_ANALIZADA <= 2'b00;
				end
			end
			
			else if (ESTADO_ACTUAL == ESTADO_MOVIENDO_HACIA_ABAJO) begin
				tableroJuego[0][0] <= 4'b1000;
				ESTADO_ACTUAL <= ESTADO_ESPERANDO_MOVIMIENTO;
			end
		end
	end
	
	// INICIO DEL CONTROL DE LOS CONTADORES.
	always @(posedge reloj) begin
		if (reinicio == 1'b1) begin
			CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_COLUMNA_ALEATORIA <= 0;
			CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_FILA_ALEATORIA <= 0;
		end
		else begin
			if (CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_COLUMNA_ALEATORIA > 22'd4000000) begin
				CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_COLUMNA_ALEATORIA <= 0;
			end
			else begin
				CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_COLUMNA_ALEATORIA <= CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_COLUMNA_ALEATORIA + 1'b1;
			end
			if (CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_FILA_ALEATORIA > 19'd400000) begin
				CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_FILA_ALEATORIA <= 0;
			end
			else begin
				CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_FILA_ALEATORIA <= CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_FILA_ALEATORIA + 1'b1;
			end
		end
	end
	// FIN DEL CONTROL DE LOS CONTADORES.

	// INICIO DEL CONTROL DE LAS POSICIONES.
	always @(posedge reloj) begin
		if (reinicio == 1'b1) begin
			POSICION_COLUMNA_ALEATORIA <= 2'd0;
			POSICION_FILA_ALEATORIA <= 2'd0;
		end
		else begin
			if (ESTADO_ACTUAL != ESTADO_GENERANDO_POSICION_ALEATORIA) begin
				if ((CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_COLUMNA_ALEATORIA >= 22'd0) && (CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_COLUMNA_ALEATORIA < 22'd1000000)) begin
					POSICION_COLUMNA_ALEATORIA <= 2'd0;
				end
				else if ((CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_COLUMNA_ALEATORIA >= 22'd1000000) && (CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_COLUMNA_ALEATORIA < 22'd2000000)) begin
					POSICION_COLUMNA_ALEATORIA <= 2'd1;
				end
				else if ((CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_COLUMNA_ALEATORIA >= 22'd2000000) && (CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_COLUMNA_ALEATORIA < 22'd3000000)) begin
					POSICION_COLUMNA_ALEATORIA <= 2'd2;
				end
				else if ((CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_COLUMNA_ALEATORIA >= 22'd3000000) && (CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_COLUMNA_ALEATORIA <= 22'd4000000)) begin
					POSICION_COLUMNA_ALEATORIA <= 2'd3;
				end
				else POSICION_COLUMNA_ALEATORIA <= 2'd3;

				if ((CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_FILA_ALEATORIA >= 19'd0) && (CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_FILA_ALEATORIA < 19'd100000)) begin
					POSICION_FILA_ALEATORIA <= 2'd0;
				end
				else if ((CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_FILA_ALEATORIA >= 19'd100000) && (CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_FILA_ALEATORIA < 19'd200000)) begin
					POSICION_FILA_ALEATORIA <= 2'd1;
				end
				else if ((CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_FILA_ALEATORIA >= 19'd200000) && (CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_FILA_ALEATORIA < 19'd300000)) begin
					POSICION_FILA_ALEATORIA <= 2'd2;
				end
				else if ((CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_FILA_ALEATORIA >= 19'd300000) && (CANTIDAD_CICLOS_RELOJ_GENERADOR_POSICION_FILA_ALEATORIA <= 19'd400000)) begin
					POSICION_FILA_ALEATORIA <= 2'd3;
				end
				else POSICION_FILA_ALEATORIA <= 2'd3; 
			end
		end
	end
	// FIN DEL CONTROL DE LAS POSICIONES.
	
	
		
endmodule 